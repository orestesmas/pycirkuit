.PS
scale=2.54
cct_init
l=elen_

# This drawing is interesting as it shows how to reuse drawing code
# This is the first stage of the filter
# Starting from left to right
In: Here
resistor(right_ 3*l/4);llabel(,R_1)
Mid: dot
resistor(right_ 3*l/4);llabel(,R_2)
dot
{
  capacitor(down_ l);rlabel(,C_1)
  GND: ground(,T,E)
}
line right_ l/2
AO: opamp(right_ 5*l/6,,,,R) with .In1 at Here
line left_ l/6 from AO.In2 then down elen_/3 then right_ elen_ then up to AO.Out
dot
line up_ 3*l/4 from AO.Out
corner
capacitor(left_ Here.x-Mid.x);rlabel(,C_2)
corner
line to Mid

# From AO's output, move slightly up and right to start the second stage
# aligned with the first
move to AO.Out
line right_ elen_/4
corner
line up_ In.y-Here.y
corner

# This is the second stage of the filter
# The code is copypasted from first stage, changing only the labels
In2: Here
resistor(right_ 3*l/4);llabel(,R_3)
Mid2: dot
resistor(right_ 3*l/4);llabel(,R_4)
dot
{
  capacitor(down_ l);rlabel(,C_3)
  GND2: ground(,T,E)
}
line right_ l/2
AO2: opamp(right_ 5*l/6,,,,R) with .In1 at Here
line left_ l/6 from AO2.In2 then down elen_/3 then right_ elen_ then up to AO2.Out
dot
line up_ 3*l/4 from AO2.Out
corner
capacitor(left_ Here.x-Mid2.x);rlabel(,C_4)
corner
line to Mid2

# The third stage is a voltage divider
move to AO2.Out
line right_ elen_/4
corner
line up_ In.y-Here.y
corner
resistor(right_ l);llabel(,R_a)
dot
{
  resistor(down_ Here.y-GND.y);rlabel(,R_b)
  ground(,T,E)
}
line right_ l/3
# Output port
dot(,,1)
# Input port (drawing it at the end avoids being overwritten by the lines starting on it)
dot(at In,,1)

.PE 
