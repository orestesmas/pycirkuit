.PS
scale=2.54
cct_init
l=elen_

In: Here
resistor(right_ 3*l/4);llabel(,R_1)
Mid: dot
resistor(right_ 3*l/4);llabel(,R_2)
dot
{
  capacitor(down_ l);rlabel(,C_1)
  GND: ground(,T,E)
}
line right_ l/2
AO: opamp(right_ 5*l/6,,,,R) with .In1 at Here
line left_ l/6 from AO.In2 then down elen_/3 then right_ elen_ then up to AO.Out
dot
#"$\,v_o(t)$" ljust
line up_ 3*l/4 from AO.Out
corner
capacitor(left_ Here.x-Mid.x);rlabel(,C_2)
corner
line to Mid
dot(at In,,1)

# Segona part
move to AO.Out
line right_ elen_/4
corner
line up_ In.y-Here.y
corner
In2: Here
resistor(right_ 3*l/4);llabel(,R_3)
Mid2: dot
resistor(right_ 3*l/4);llabel(,R_4)
dot
{
  capacitor(down_ l);rlabel(,C_3)
  GND2: ground(,T,E)
}
line right_ l/2
AO2: opamp(right_ 5*l/6,,,,R) with .In1 at Here
line left_ l/6 from AO2.In2 then down elen_/3 then right_ elen_ then up to AO2.Out
dot
line up_ 3*l/4 from AO2.Out
corner
capacitor(left_ Here.x-Mid2.x);rlabel(,C_4)
corner
line to Mid2

# Tercera etapa
move to AO2.Out
line right_ elen_/4
corner
line up_ In.y-Here.y
corner
resistor(right_ l);llabel(,R_a)
dot
{
  resistor(down_ Here.y-GND.y);rlabel(,R_b)
  ground(,T,E)
}
line right_ l/3
dot(,,1)

.PE 
